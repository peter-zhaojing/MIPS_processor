module MIPS150(
	input 	clk, rst,
	input		FPGA_SERIAL_RX,
	output	FPGA_SERIAL_TX
);

// Use this as the top-level module for your CPU. You
// will likely want to break control and datapath out
// into separate modules that you instantiate here.

//declare signals for connection
wire	[31:0]	Instr;
wire	[3:0]		ALUControl;
wire				RegWrite;
wire	[2:0]		Mask;
wire  [1:0]		MemWrite;
wire				MemtoReg;
wire				LUItoReg;
wire				SignOrZero;
wire				ALUSrc;
wire				RegDst;
wire				VarOrShamt;
wire	[2:0]		BranchCtrl;
wire				Jump;
wire				JAL;
wire				JLink;
wire				JumpReg;

//instantiate datapath
MIPS150_datapath mips_datapath(
	.clk			(clk),
	.rst			(rst),
	.Instr		(Instr),
	.ALUControl	(ALUControl),
	.RegWrite	(RegWrite),
	.Mask			(Mask),
	.MemWrite	(MemWrite),
	.MemtoReg	(MemtoReg),
	.LUItoReg	(LUItoReg),
	.SignOrZero	(SignOrZero),
	.ALUSrc		(ALUSrc),
	.RegDst		(RegDst),
	.VarOrShamt	(VarOrShamt),
	.BranchCtrl	(BranchCtrl),
	.Jump			(Jump),
	.JAL			(JAL),
	.JLink		(JLink),
	.JumpReg		(JumpReg)
);


//instantiate control unit
MIPS150_control mips_control(
	 .Instr			(Instr),
	 .ALUControl	(ALUControl),
	 .RegWrite		(RegWrite),
	 .Mask			(Mask),
	 .MemWrite		(MemWrite),
	 .MemtoReg		(MemtoReg),
	 .LUItoReg		(LUItoReg),
	 .SignOrZero	(SignOrZero),
	 .ALUSrc			(ALUSrc),
	 .RegDst			(RegDst),
	 .VarOrShamt	(VarOrShamt),
	 .BranchCtrl	(BranchCtrl),
	 .Jump			(Jump),
	 .JAL				(JAL),
	 .JLink			(JLink),
	 .JumpReg		(JumpReg)
);

endmodule
